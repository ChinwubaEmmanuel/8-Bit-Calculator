module calc_out(
input [7:0] A,
input LoadOU, clock,
//input clock, reset, OnOff,
output a1,b1,c1,d1,e1,f1,g1,a2,b2,c2,d2,e2,f2,g2,a3,b3,c3,d3,e3,f3,g3,a4,b4,c4,d4,e4,f4,g4
);
//wire clk;
//wire [8:0] testpatt;
reg [3:0] SB;
wire [7:0] S;
wire [3:0] ONES, TENS;
wire [1:0] HUNDREDS;
/*
OneHertzClock
(
	.clock(clock) ,	// input  clock_sig
	.reset(reset) ,	// input  reset_sig
	.OnOff(OnOff) ,	// input  OnOff_sig
	.FinalOneHertz(clk) 	// output  FinalOneHertz_sig
);

divideXn #(10'd256, 4'd9) div8
(
	.CLK(clk) ,	// input  CLK_sig
	.CLEAR(reset) ,	// input  CLEAR_sig
	.COUNT(testpatt) ,	// output [M-1:0] COUNT_sig
	.OUT(out) 	// output  OUT_sig
);

MUX_reg
(
	.y(D) ,	// output [7:0] y_sig
	.a(A) ,	// input [7:0] a_sig
	.load(LoadOU) ,	// input  load_sig
	.clear(reset) 	// input  clear_sig
);
NbitOU NbitOU_inst1
(
	.D(A) ,	// input [N-1:0] D_sig
	.Load(LoadOU) ,	// input  Load_sig
	.clr(reset) ,	// input  clr_sig
	.clock(clock) ,	// input  clock_sig
	.Q(D) 	// output [N-1:0] Q_sig
); */
calc_out_unit signmag
(
	.a(A) ,	// input [7:0] a_sig
	.s(S) 	// output [7:0] s_sig
);
binary2bcd
(
	.A({1'b0,S[6:0]}) ,	// input [7:0] A_sig
	.ONES(ONES) ,	// output [3:0] ONES_sig
	.TENS(TENS) ,	// output [3:0] TENS_sig
	.HUNDREDS(HUNDREDS) 	// output [1:0] HUNDREDS_sig
);

binary2seven
(
	.w(ONES[3]) ,	// input  w_sig
	.x(ONES[2]) ,	// input  x_sig
	.y(ONES[1]) ,	// input  y_sig
	.z(ONES[0]) ,	// input  z_sig
	.a(a1) ,	// output  a_sig
	.b(b1) ,	// output  b_sig
	.c(c1) ,	// output  c_sig
	.d(d1) ,	// output  d_sig
	.e(e1) ,	// output  e_sig
	.f(f1) ,	// output  f_sig
	.g(g1) 	// output  g_sig
);

binary2seven
(
	.w(TENS[3]) ,	// input  w_sig
	.x(TENS[2]) ,	// input  x_sig
	.y(TENS[1]) ,	// input  y_sig
	.z(TENS[0]) ,	// input  z_sig
	.a(a2) ,	// output  a_sig
	.b(b2) ,	// output  b_sig
	.c(c2) ,	// output  c_sig
	.d(d2) ,	// output  d_sig
	.e(e2) ,	// output  e_sig
	.f(f2) ,	// output  f_sig
	.g(g2) 	// output  g_sig
);
binary2seven
(
	.w(1'b0) ,	// input  w_sig
	.x(1'b0) ,	// input  x_sig
	.y(HUNDREDS[1]) ,	// input  y_sig
	.z(HUNDREDS[0]) ,	// input  z_sig
	.a(a3) ,	// output  a_sig
	.b(b3) ,	// output  b_sig
	.c(c3) ,	// output  c_sig
	.d(d3) ,	// output  d_sig
	.e(e3) ,	// output  e_sig
	.f(f3) ,	// output  f_sig
	.g(g3) 	// output  g_sig
);

always @ (A) begin
	if(A[7] == 1) begin
		SB[0] = 1;
		SB[1] = 1;
		SB[2] = 1;
		SB[3] = 1;
end	else begin
		SB[0] = 0;
		SB[1] = 1;
		SB[2] = 1;
		SB[3] = 1;
	end
end

binary2seven
(
	.w(SB[3]) ,	// input  w_sig
	.x(SB[2]) ,	// input  x_sig
	.y(SB[1]) ,	// input  y_sig
	.z(SB[0]) ,	// input  z_sig
	.a(a4) ,	// output  a_sig
	.b(b4) ,	// output  b_sig
	.c(c4) ,	// output  c_sig
	.d(d4) ,	// output  d_sig
	.e(e4) ,	// output  e_sig
	.f(f4) ,	// output  f_sig
	.g(g4) 	// output  g_sig
);
endmodule